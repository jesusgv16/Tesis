library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity SIGMAGRANDE1 is
	 port(
		 EX : in  STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SF : out STD_LOGIC_VECTOR(31 DOWNTO 0)
	     );
end SIGMAGRANDE1;
 
architecture SIGMAGRANDE1 of SIGMAGRANDE1 is
COMPONENT XOR2TO1_32BIT is
	 port(
		 EX1 : in STD_LOGIC_VECTOR(31 downto 0);
		 EX2 : in STD_LOGIC_VECTOR(31 downto 0);
		 SX : out STD_LOGIC_VECTOR(31 downto 0)
	     );
end COMPONENT;		   
SIGNAL SX1: STD_LOGIC_VECTOR (31 DOWNTO 0);
begin	   
	XOR1: XOR2TO1_32BIT PORT MAP (
		EX1(31 DOWNTO 26)=>EX( 5 DOWNTO 0),
		EX1(25 DOWNTO  0)=>EX(31 DOWNTO 6),
		EX2(31 DOWNTO 21)=>EX(10 DOWNTO 0),
		EX2(20 DOWNTO  0)=>EX(31 DOWNTO 11),
		SX =>SX1
		);
	XOR2: XOR2TO1_32BIT PORT MAP (
		EX1(31 DOWNTO  7)=>EX(24 DOWNTO 0),
		EX1( 6 DOWNTO  0)=>EX(31 DOWNTO 25),
		EX2=>SX1,
		SX =>SF
		);
end SIGMAGRANDE1;