---------------------------------------------------------------------------------------------------
--
-- Title       : REGTEMP_128BIT
-- Design      : AES_IAB27
-- Author      : IAB27
-- Company     : INAOE
--
---------------------------------------------------------------------------------------------------
--
-- File        : REGTEMP_128BIT.vhd
-- Generated   : Mon Jan 12 10:28:57 2004
-- From        : TLAX
-- By          : AZTEC Ver. 1.0
--
---------------------------------------------------------------------------------------------------
--
-- Description : 
--
---------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity REGTEMP_128BIT is
	 port(
		 ERD : in STD_LOGIC_VECTOR(127 downto 0);
		 ERW : in STD_LOGIC;
		 CLK : in STD_LOGIC;
		 RST : in STD_LOGIC;
		 SRQ : out STD_LOGIC_VECTOR(127 downto 0)
	     );
end REGTEMP_128BIT;

architecture REGTEMP_128BIT of REGTEMP_128BIT is
	component REGTEMP_1BIT is
	 port(
		 ERD : in STD_LOGIC;
		 ERW : in STD_LOGIC;
		 CLK : in STD_LOGIC;
		 RST : in STD_LOGIC;
		 SRQ : out STD_LOGIC
	     );
	end component;
begin
	R000: REGTEMP_1BIT PORT MAP (ERD(  0),ERW,CLK,RST,SRQ(  0));
	R001: REGTEMP_1BIT PORT MAP (ERD(  1),ERW,CLK,RST,SRQ(  1));
	R002: REGTEMP_1BIT PORT MAP (ERD(  2),ERW,CLK,RST,SRQ(  2));
	R003: REGTEMP_1BIT PORT MAP (ERD(  3),ERW,CLK,RST,SRQ(  3));
	R004: REGTEMP_1BIT PORT MAP (ERD(  4),ERW,CLK,RST,SRQ(  4));
	R005: REGTEMP_1BIT PORT MAP (ERD(  5),ERW,CLK,RST,SRQ(  5));
	R006: REGTEMP_1BIT PORT MAP (ERD(  6),ERW,CLK,RST,SRQ(  6));
	R007: REGTEMP_1BIT PORT MAP (ERD(  7),ERW,CLK,RST,SRQ(  7));
	R008: REGTEMP_1BIT PORT MAP (ERD(  8),ERW,CLK,RST,SRQ(  8));
	R009: REGTEMP_1BIT PORT MAP (ERD(  9),ERW,CLK,RST,SRQ(  9));
	R010: REGTEMP_1BIT PORT MAP (ERD( 10),ERW,CLK,RST,SRQ( 10));
	R011: REGTEMP_1BIT PORT MAP (ERD( 11),ERW,CLK,RST,SRQ( 11));
	R012: REGTEMP_1BIT PORT MAP (ERD( 12),ERW,CLK,RST,SRQ( 12));
	R013: REGTEMP_1BIT PORT MAP (ERD( 13),ERW,CLK,RST,SRQ( 13));
	R014: REGTEMP_1BIT PORT MAP (ERD( 14),ERW,CLK,RST,SRQ( 14));
	R015: REGTEMP_1BIT PORT MAP (ERD( 15),ERW,CLK,RST,SRQ( 15));
	R016: REGTEMP_1BIT PORT MAP (ERD( 16),ERW,CLK,RST,SRQ( 16));
	R017: REGTEMP_1BIT PORT MAP (ERD( 17),ERW,CLK,RST,SRQ( 17));
	R018: REGTEMP_1BIT PORT MAP (ERD( 18),ERW,CLK,RST,SRQ( 18));
	R019: REGTEMP_1BIT PORT MAP (ERD( 19),ERW,CLK,RST,SRQ( 19));
	R020: REGTEMP_1BIT PORT MAP (ERD( 20),ERW,CLK,RST,SRQ( 20));
	R021: REGTEMP_1BIT PORT MAP (ERD( 21),ERW,CLK,RST,SRQ( 21));
	R022: REGTEMP_1BIT PORT MAP (ERD( 22),ERW,CLK,RST,SRQ( 22));
	R023: REGTEMP_1BIT PORT MAP (ERD( 23),ERW,CLK,RST,SRQ( 23));
	R024: REGTEMP_1BIT PORT MAP (ERD( 24),ERW,CLK,RST,SRQ( 24));
	R025: REGTEMP_1BIT PORT MAP (ERD( 25),ERW,CLK,RST,SRQ( 25));
	R026: REGTEMP_1BIT PORT MAP (ERD( 26),ERW,CLK,RST,SRQ( 26));
	R027: REGTEMP_1BIT PORT MAP (ERD( 27),ERW,CLK,RST,SRQ( 27));
	R028: REGTEMP_1BIT PORT MAP (ERD( 28),ERW,CLK,RST,SRQ( 28));
	R029: REGTEMP_1BIT PORT MAP (ERD( 29),ERW,CLK,RST,SRQ( 29));
	R030: REGTEMP_1BIT PORT MAP (ERD( 30),ERW,CLK,RST,SRQ( 30));
	R031: REGTEMP_1BIT PORT MAP (ERD( 31),ERW,CLK,RST,SRQ( 31));
	R032: REGTEMP_1BIT PORT MAP (ERD( 32),ERW,CLK,RST,SRQ( 32));
	R033: REGTEMP_1BIT PORT MAP (ERD( 33),ERW,CLK,RST,SRQ( 33));
	R034: REGTEMP_1BIT PORT MAP (ERD( 34),ERW,CLK,RST,SRQ( 34));
	R035: REGTEMP_1BIT PORT MAP (ERD( 35),ERW,CLK,RST,SRQ( 35));
	R036: REGTEMP_1BIT PORT MAP (ERD( 36),ERW,CLK,RST,SRQ( 36));
	R037: REGTEMP_1BIT PORT MAP (ERD( 37),ERW,CLK,RST,SRQ( 37));
	R038: REGTEMP_1BIT PORT MAP (ERD( 38),ERW,CLK,RST,SRQ( 38));
	R039: REGTEMP_1BIT PORT MAP (ERD( 39),ERW,CLK,RST,SRQ( 39));
	R040: REGTEMP_1BIT PORT MAP (ERD( 40),ERW,CLK,RST,SRQ( 40));
	R041: REGTEMP_1BIT PORT MAP (ERD( 41),ERW,CLK,RST,SRQ( 41));
	R042: REGTEMP_1BIT PORT MAP (ERD( 42),ERW,CLK,RST,SRQ( 42));
	R043: REGTEMP_1BIT PORT MAP (ERD( 43),ERW,CLK,RST,SRQ( 43));
	R044: REGTEMP_1BIT PORT MAP (ERD( 44),ERW,CLK,RST,SRQ( 44));
	R045: REGTEMP_1BIT PORT MAP (ERD( 45),ERW,CLK,RST,SRQ( 45));
	R046: REGTEMP_1BIT PORT MAP (ERD( 46),ERW,CLK,RST,SRQ( 46));
	R047: REGTEMP_1BIT PORT MAP (ERD( 47),ERW,CLK,RST,SRQ( 47));
	R048: REGTEMP_1BIT PORT MAP (ERD( 48),ERW,CLK,RST,SRQ( 48));
	R049: REGTEMP_1BIT PORT MAP (ERD( 49),ERW,CLK,RST,SRQ( 49));
	R050: REGTEMP_1BIT PORT MAP (ERD( 50),ERW,CLK,RST,SRQ( 50));
	R051: REGTEMP_1BIT PORT MAP (ERD( 51),ERW,CLK,RST,SRQ( 51));
	R052: REGTEMP_1BIT PORT MAP (ERD( 52),ERW,CLK,RST,SRQ( 52));
	R053: REGTEMP_1BIT PORT MAP (ERD( 53),ERW,CLK,RST,SRQ( 53));
	R054: REGTEMP_1BIT PORT MAP (ERD( 54),ERW,CLK,RST,SRQ( 54));
	R055: REGTEMP_1BIT PORT MAP (ERD( 55),ERW,CLK,RST,SRQ( 55));
	R056: REGTEMP_1BIT PORT MAP (ERD( 56),ERW,CLK,RST,SRQ( 56));
	R057: REGTEMP_1BIT PORT MAP (ERD( 57),ERW,CLK,RST,SRQ( 57));
	R058: REGTEMP_1BIT PORT MAP (ERD( 58),ERW,CLK,RST,SRQ( 58));
	R059: REGTEMP_1BIT PORT MAP (ERD( 59),ERW,CLK,RST,SRQ( 59));
	R060: REGTEMP_1BIT PORT MAP (ERD( 60),ERW,CLK,RST,SRQ( 60));
	R061: REGTEMP_1BIT PORT MAP (ERD( 61),ERW,CLK,RST,SRQ( 61));
	R062: REGTEMP_1BIT PORT MAP (ERD( 62),ERW,CLK,RST,SRQ( 62));
	R063: REGTEMP_1BIT PORT MAP (ERD( 63),ERW,CLK,RST,SRQ( 63));
	R064: REGTEMP_1BIT PORT MAP (ERD( 64),ERW,CLK,RST,SRQ( 64));
	R065: REGTEMP_1BIT PORT MAP (ERD( 65),ERW,CLK,RST,SRQ( 65));
	R066: REGTEMP_1BIT PORT MAP (ERD( 66),ERW,CLK,RST,SRQ( 66));
	R067: REGTEMP_1BIT PORT MAP (ERD( 67),ERW,CLK,RST,SRQ( 67));
	R068: REGTEMP_1BIT PORT MAP (ERD( 68),ERW,CLK,RST,SRQ( 68));
	R069: REGTEMP_1BIT PORT MAP (ERD( 69),ERW,CLK,RST,SRQ( 69));
	R070: REGTEMP_1BIT PORT MAP (ERD( 70),ERW,CLK,RST,SRQ( 70));
	R071: REGTEMP_1BIT PORT MAP (ERD( 71),ERW,CLK,RST,SRQ( 71));
	R072: REGTEMP_1BIT PORT MAP (ERD( 72),ERW,CLK,RST,SRQ( 72));
	R073: REGTEMP_1BIT PORT MAP (ERD( 73),ERW,CLK,RST,SRQ( 73));
	R074: REGTEMP_1BIT PORT MAP (ERD( 74),ERW,CLK,RST,SRQ( 74));
	R075: REGTEMP_1BIT PORT MAP (ERD( 75),ERW,CLK,RST,SRQ( 75));
	R076: REGTEMP_1BIT PORT MAP (ERD( 76),ERW,CLK,RST,SRQ( 76));
	R077: REGTEMP_1BIT PORT MAP (ERD( 77),ERW,CLK,RST,SRQ( 77));
	R078: REGTEMP_1BIT PORT MAP (ERD( 78),ERW,CLK,RST,SRQ( 78));
	R079: REGTEMP_1BIT PORT MAP (ERD( 79),ERW,CLK,RST,SRQ( 79));
	R080: REGTEMP_1BIT PORT MAP (ERD( 80),ERW,CLK,RST,SRQ( 80));
	R081: REGTEMP_1BIT PORT MAP (ERD( 81),ERW,CLK,RST,SRQ( 81));
	R082: REGTEMP_1BIT PORT MAP (ERD( 82),ERW,CLK,RST,SRQ( 82));
	R083: REGTEMP_1BIT PORT MAP (ERD( 83),ERW,CLK,RST,SRQ( 83));
	R084: REGTEMP_1BIT PORT MAP (ERD( 84),ERW,CLK,RST,SRQ( 84));
	R085: REGTEMP_1BIT PORT MAP (ERD( 85),ERW,CLK,RST,SRQ( 85));
	R086: REGTEMP_1BIT PORT MAP (ERD( 86),ERW,CLK,RST,SRQ( 86));
	R087: REGTEMP_1BIT PORT MAP (ERD( 87),ERW,CLK,RST,SRQ( 87));
	R088: REGTEMP_1BIT PORT MAP (ERD( 88),ERW,CLK,RST,SRQ( 88));
	R089: REGTEMP_1BIT PORT MAP (ERD( 89),ERW,CLK,RST,SRQ( 89));
	R090: REGTEMP_1BIT PORT MAP (ERD( 90),ERW,CLK,RST,SRQ( 90));
	R091: REGTEMP_1BIT PORT MAP (ERD( 91),ERW,CLK,RST,SRQ( 91));
	R092: REGTEMP_1BIT PORT MAP (ERD( 92),ERW,CLK,RST,SRQ( 92));
	R093: REGTEMP_1BIT PORT MAP (ERD( 93),ERW,CLK,RST,SRQ( 93));
	R094: REGTEMP_1BIT PORT MAP (ERD( 94),ERW,CLK,RST,SRQ( 94));
	R095: REGTEMP_1BIT PORT MAP (ERD( 95),ERW,CLK,RST,SRQ( 95));
	R096: REGTEMP_1BIT PORT MAP (ERD( 96),ERW,CLK,RST,SRQ( 96));
	R097: REGTEMP_1BIT PORT MAP (ERD( 97),ERW,CLK,RST,SRQ( 97));
	R098: REGTEMP_1BIT PORT MAP (ERD( 98),ERW,CLK,RST,SRQ( 98));
	R099: REGTEMP_1BIT PORT MAP (ERD( 99),ERW,CLK,RST,SRQ( 99));
	R100: REGTEMP_1BIT PORT MAP (ERD(100),ERW,CLK,RST,SRQ(100));
	R101: REGTEMP_1BIT PORT MAP (ERD(101),ERW,CLK,RST,SRQ(101));
	R102: REGTEMP_1BIT PORT MAP (ERD(102),ERW,CLK,RST,SRQ(102));
	R103: REGTEMP_1BIT PORT MAP (ERD(103),ERW,CLK,RST,SRQ(103));
	R104: REGTEMP_1BIT PORT MAP (ERD(104),ERW,CLK,RST,SRQ(104));
	R105: REGTEMP_1BIT PORT MAP (ERD(105),ERW,CLK,RST,SRQ(105));
	R106: REGTEMP_1BIT PORT MAP (ERD(106),ERW,CLK,RST,SRQ(106));
	R107: REGTEMP_1BIT PORT MAP (ERD(107),ERW,CLK,RST,SRQ(107));
	R108: REGTEMP_1BIT PORT MAP (ERD(108),ERW,CLK,RST,SRQ(108));
	R109: REGTEMP_1BIT PORT MAP (ERD(109),ERW,CLK,RST,SRQ(109));
	R110: REGTEMP_1BIT PORT MAP (ERD(110),ERW,CLK,RST,SRQ(110));
	R111: REGTEMP_1BIT PORT MAP (ERD(111),ERW,CLK,RST,SRQ(111));
	R112: REGTEMP_1BIT PORT MAP (ERD(112),ERW,CLK,RST,SRQ(112));
	R113: REGTEMP_1BIT PORT MAP (ERD(113),ERW,CLK,RST,SRQ(113));
	R114: REGTEMP_1BIT PORT MAP (ERD(114),ERW,CLK,RST,SRQ(114));
	R115: REGTEMP_1BIT PORT MAP (ERD(115),ERW,CLK,RST,SRQ(115));
	R116: REGTEMP_1BIT PORT MAP (ERD(116),ERW,CLK,RST,SRQ(116));
	R117: REGTEMP_1BIT PORT MAP (ERD(117),ERW,CLK,RST,SRQ(117));
	R118: REGTEMP_1BIT PORT MAP (ERD(118),ERW,CLK,RST,SRQ(118));
	R119: REGTEMP_1BIT PORT MAP (ERD(119),ERW,CLK,RST,SRQ(119));
	R120: REGTEMP_1BIT PORT MAP (ERD(120),ERW,CLK,RST,SRQ(120));
	R121: REGTEMP_1BIT PORT MAP (ERD(121),ERW,CLK,RST,SRQ(121));
	R122: REGTEMP_1BIT PORT MAP (ERD(122),ERW,CLK,RST,SRQ(122));
	R123: REGTEMP_1BIT PORT MAP (ERD(123),ERW,CLK,RST,SRQ(123));
	R124: REGTEMP_1BIT PORT MAP (ERD(124),ERW,CLK,RST,SRQ(124));
	R125: REGTEMP_1BIT PORT MAP (ERD(125),ERW,CLK,RST,SRQ(125));
	R126: REGTEMP_1BIT PORT MAP (ERD(126),ERW,CLK,RST,SRQ(126));
	R127: REGTEMP_1BIT PORT MAP (ERD(127),ERW,CLK,RST,SRQ(127));
end REGTEMP_128BIT;
