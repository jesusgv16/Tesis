---------------------------------------------------------------------------------------------------
--
-- Title       : MUX2TO1_128BIT
-- Design      : MD5_IAB27_B
-- Author      : IAB27
-- Company     : Home
--
---------------------------------------------------------------------------------------------------
--
-- File        : MUX2TO1_128BIT.vhd
-- Generated   : Tue Feb 24 20:54:41 2004
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.20
--
---------------------------------------------------------------------------------------------------
--
-- Description : 
--
---------------------------------------------------------------------------------------------------
 
library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity MUX2TO1_128BIT is
	 port(
		 EM1 : in STD_LOGIC_VECTOR(127 downto 0);
		 EM2 : in STD_LOGIC_VECTOR(127 downto 0);
		 EMS : in STD_LOGIC;
		 SM : out STD_LOGIC_VECTOR(127 downto 0)
	     );
end MUX2TO1_128BIT;
 
architecture MUX2TO1_128BIT of MUX2TO1_128BIT is
component MUX2TO1_1BIT is
	 port(
		 EM1 : in STD_LOGIC;
		 EM2 : in STD_LOGIC;
		 EMS : in STD_LOGIC;
		 SM : out STD_LOGIC
	     );
	end component;
begin
	M000: MUX2TO1_1BIT PORT MAP (EM1(  0),EM2(  0),EMS,SM(  0));
	M001: MUX2TO1_1BIT PORT MAP (EM1(  1),EM2(  1),EMS,SM(  1));
	M002: MUX2TO1_1BIT PORT MAP (EM1(  2),EM2(  2),EMS,SM(  2));
	M003: MUX2TO1_1BIT PORT MAP (EM1(  3),EM2(  3),EMS,SM(  3));
	M004: MUX2TO1_1BIT PORT MAP (EM1(  4),EM2(  4),EMS,SM(  4));
	M005: MUX2TO1_1BIT PORT MAP (EM1(  5),EM2(  5),EMS,SM(  5));
	M006: MUX2TO1_1BIT PORT MAP (EM1(  6),EM2(  6),EMS,SM(  6));
	M007: MUX2TO1_1BIT PORT MAP (EM1(  7),EM2(  7),EMS,SM(  7));
	M008: MUX2TO1_1BIT PORT MAP (EM1(  8),EM2(  8),EMS,SM(  8));
	M009: MUX2TO1_1BIT PORT MAP (EM1(  9),EM2(  9),EMS,SM(  9));
	M010: MUX2TO1_1BIT PORT MAP (EM1( 10),EM2( 10),EMS,SM( 10));
	M011: MUX2TO1_1BIT PORT MAP (EM1( 11),EM2( 11),EMS,SM( 11));
	M012: MUX2TO1_1BIT PORT MAP (EM1( 12),EM2( 12),EMS,SM( 12));
	M013: MUX2TO1_1BIT PORT MAP (EM1( 13),EM2( 13),EMS,SM( 13));
	M014: MUX2TO1_1BIT PORT MAP (EM1( 14),EM2( 14),EMS,SM( 14));
	M015: MUX2TO1_1BIT PORT MAP (EM1( 15),EM2( 15),EMS,SM( 15));
	M016: MUX2TO1_1BIT PORT MAP (EM1( 16),EM2( 16),EMS,SM( 16));
	M017: MUX2TO1_1BIT PORT MAP (EM1( 17),EM2( 17),EMS,SM( 17));
	M018: MUX2TO1_1BIT PORT MAP (EM1( 18),EM2( 18),EMS,SM( 18));
	M019: MUX2TO1_1BIT PORT MAP (EM1( 19),EM2( 19),EMS,SM( 19));
	M020: MUX2TO1_1BIT PORT MAP (EM1( 20),EM2( 20),EMS,SM( 20));
	M021: MUX2TO1_1BIT PORT MAP (EM1( 21),EM2( 21),EMS,SM( 21));
	M022: MUX2TO1_1BIT PORT MAP (EM1( 22),EM2( 22),EMS,SM( 22));
	M023: MUX2TO1_1BIT PORT MAP (EM1( 23),EM2( 23),EMS,SM( 23));
	M024: MUX2TO1_1BIT PORT MAP (EM1( 24),EM2( 24),EMS,SM( 24));
	M025: MUX2TO1_1BIT PORT MAP (EM1( 25),EM2( 25),EMS,SM( 25));
	M026: MUX2TO1_1BIT PORT MAP (EM1( 26),EM2( 26),EMS,SM( 26));
	M027: MUX2TO1_1BIT PORT MAP (EM1( 27),EM2( 27),EMS,SM( 27));
	M028: MUX2TO1_1BIT PORT MAP (EM1( 28),EM2( 28),EMS,SM( 28));
	M029: MUX2TO1_1BIT PORT MAP (EM1( 29),EM2( 29),EMS,SM( 29));
	M030: MUX2TO1_1BIT PORT MAP (EM1( 30),EM2( 30),EMS,SM( 30));
	M031: MUX2TO1_1BIT PORT MAP (EM1( 31),EM2( 31),EMS,SM( 31));
	M032: MUX2TO1_1BIT PORT MAP (EM1( 32),EM2( 32),EMS,SM( 32));
	M033: MUX2TO1_1BIT PORT MAP (EM1( 33),EM2( 33),EMS,SM( 33));
	M034: MUX2TO1_1BIT PORT MAP (EM1( 34),EM2( 34),EMS,SM( 34));
	M035: MUX2TO1_1BIT PORT MAP (EM1( 35),EM2( 35),EMS,SM( 35));
	M036: MUX2TO1_1BIT PORT MAP (EM1( 36),EM2( 36),EMS,SM( 36));
	M037: MUX2TO1_1BIT PORT MAP (EM1( 37),EM2( 37),EMS,SM( 37));
	M038: MUX2TO1_1BIT PORT MAP (EM1( 38),EM2( 38),EMS,SM( 38));
	M039: MUX2TO1_1BIT PORT MAP (EM1( 39),EM2( 39),EMS,SM( 39));
	M040: MUX2TO1_1BIT PORT MAP (EM1( 40),EM2( 40),EMS,SM( 40));
	M041: MUX2TO1_1BIT PORT MAP (EM1( 41),EM2( 41),EMS,SM( 41));
	M042: MUX2TO1_1BIT PORT MAP (EM1( 42),EM2( 42),EMS,SM( 42));
	M043: MUX2TO1_1BIT PORT MAP (EM1( 43),EM2( 43),EMS,SM( 43));
	M044: MUX2TO1_1BIT PORT MAP (EM1( 44),EM2( 44),EMS,SM( 44));
	M045: MUX2TO1_1BIT PORT MAP (EM1( 45),EM2( 45),EMS,SM( 45));
	M046: MUX2TO1_1BIT PORT MAP (EM1( 46),EM2( 46),EMS,SM( 46));
	M047: MUX2TO1_1BIT PORT MAP (EM1( 47),EM2( 47),EMS,SM( 47));
	M048: MUX2TO1_1BIT PORT MAP (EM1( 48),EM2( 48),EMS,SM( 48));
	M049: MUX2TO1_1BIT PORT MAP (EM1( 49),EM2( 49),EMS,SM( 49));
	M050: MUX2TO1_1BIT PORT MAP (EM1( 50),EM2( 50),EMS,SM( 50));
	M051: MUX2TO1_1BIT PORT MAP (EM1( 51),EM2( 51),EMS,SM( 51));
	M052: MUX2TO1_1BIT PORT MAP (EM1( 52),EM2( 52),EMS,SM( 52));
	M053: MUX2TO1_1BIT PORT MAP (EM1( 53),EM2( 53),EMS,SM( 53));
	M054: MUX2TO1_1BIT PORT MAP (EM1( 54),EM2( 54),EMS,SM( 54));
	M055: MUX2TO1_1BIT PORT MAP (EM1( 55),EM2( 55),EMS,SM( 55));
	M056: MUX2TO1_1BIT PORT MAP (EM1( 56),EM2( 56),EMS,SM( 56));
	M057: MUX2TO1_1BIT PORT MAP (EM1( 57),EM2( 57),EMS,SM( 57));
	M058: MUX2TO1_1BIT PORT MAP (EM1( 58),EM2( 58),EMS,SM( 58));
	M059: MUX2TO1_1BIT PORT MAP (EM1( 59),EM2( 59),EMS,SM( 59));
	M060: MUX2TO1_1BIT PORT MAP (EM1( 60),EM2( 60),EMS,SM( 60));
	M061: MUX2TO1_1BIT PORT MAP (EM1( 61),EM2( 61),EMS,SM( 61));
	M062: MUX2TO1_1BIT PORT MAP (EM1( 62),EM2( 62),EMS,SM( 62));
	M063: MUX2TO1_1BIT PORT MAP (EM1( 63),EM2( 63),EMS,SM( 63));
	M064: MUX2TO1_1BIT PORT MAP (EM1( 64),EM2( 64),EMS,SM( 64));
	M065: MUX2TO1_1BIT PORT MAP (EM1( 65),EM2( 65),EMS,SM( 65));
	M066: MUX2TO1_1BIT PORT MAP (EM1( 66),EM2( 66),EMS,SM( 66));
	M067: MUX2TO1_1BIT PORT MAP (EM1( 67),EM2( 67),EMS,SM( 67));
	M068: MUX2TO1_1BIT PORT MAP (EM1( 68),EM2( 68),EMS,SM( 68));
	M069: MUX2TO1_1BIT PORT MAP (EM1( 69),EM2( 69),EMS,SM( 69));
	M070: MUX2TO1_1BIT PORT MAP (EM1( 70),EM2( 70),EMS,SM( 70));
	M071: MUX2TO1_1BIT PORT MAP (EM1( 71),EM2( 71),EMS,SM( 71));
	M072: MUX2TO1_1BIT PORT MAP (EM1( 72),EM2( 72),EMS,SM( 72));
	M073: MUX2TO1_1BIT PORT MAP (EM1( 73),EM2( 73),EMS,SM( 73));
	M074: MUX2TO1_1BIT PORT MAP (EM1( 74),EM2( 74),EMS,SM( 74));
	M075: MUX2TO1_1BIT PORT MAP (EM1( 75),EM2( 75),EMS,SM( 75));
	M076: MUX2TO1_1BIT PORT MAP (EM1( 76),EM2( 76),EMS,SM( 76));
	M077: MUX2TO1_1BIT PORT MAP (EM1( 77),EM2( 77),EMS,SM( 77));
	M078: MUX2TO1_1BIT PORT MAP (EM1( 78),EM2( 78),EMS,SM( 78));
	M079: MUX2TO1_1BIT PORT MAP (EM1( 79),EM2( 79),EMS,SM( 79));
	M080: MUX2TO1_1BIT PORT MAP (EM1( 80),EM2( 80),EMS,SM( 80));
	M081: MUX2TO1_1BIT PORT MAP (EM1( 81),EM2( 81),EMS,SM( 81));
	M082: MUX2TO1_1BIT PORT MAP (EM1( 82),EM2( 82),EMS,SM( 82));
	M083: MUX2TO1_1BIT PORT MAP (EM1( 83),EM2( 83),EMS,SM( 83));
	M084: MUX2TO1_1BIT PORT MAP (EM1( 84),EM2( 84),EMS,SM( 84));
	M085: MUX2TO1_1BIT PORT MAP (EM1( 85),EM2( 85),EMS,SM( 85));
	M086: MUX2TO1_1BIT PORT MAP (EM1( 86),EM2( 86),EMS,SM( 86));
	M087: MUX2TO1_1BIT PORT MAP (EM1( 87),EM2( 87),EMS,SM( 87));
	M088: MUX2TO1_1BIT PORT MAP (EM1( 88),EM2( 88),EMS,SM( 88));
	M089: MUX2TO1_1BIT PORT MAP (EM1( 89),EM2( 89),EMS,SM( 89));
	M090: MUX2TO1_1BIT PORT MAP (EM1( 90),EM2( 90),EMS,SM( 90));
	M091: MUX2TO1_1BIT PORT MAP (EM1( 91),EM2( 91),EMS,SM( 91));
	M092: MUX2TO1_1BIT PORT MAP (EM1( 92),EM2( 92),EMS,SM( 92));
	M093: MUX2TO1_1BIT PORT MAP (EM1( 93),EM2( 93),EMS,SM( 93));
	M094: MUX2TO1_1BIT PORT MAP (EM1( 94),EM2( 94),EMS,SM( 94));
	M095: MUX2TO1_1BIT PORT MAP (EM1( 95),EM2( 95),EMS,SM( 95));
	M096: MUX2TO1_1BIT PORT MAP (EM1( 96),EM2( 96),EMS,SM( 96));
	M097: MUX2TO1_1BIT PORT MAP (EM1( 97),EM2( 97),EMS,SM( 97));
	M098: MUX2TO1_1BIT PORT MAP (EM1( 98),EM2( 98),EMS,SM( 98));
	M099: MUX2TO1_1BIT PORT MAP (EM1( 99),EM2( 99),EMS,SM( 99));
	M100: MUX2TO1_1BIT PORT MAP (EM1(100),EM2(100),EMS,SM(100));
	M101: MUX2TO1_1BIT PORT MAP (EM1(101),EM2(101),EMS,SM(101));
	M102: MUX2TO1_1BIT PORT MAP (EM1(102),EM2(102),EMS,SM(102));
	M103: MUX2TO1_1BIT PORT MAP (EM1(103),EM2(103),EMS,SM(103));
	M104: MUX2TO1_1BIT PORT MAP (EM1(104),EM2(104),EMS,SM(104));
	M105: MUX2TO1_1BIT PORT MAP (EM1(105),EM2(105),EMS,SM(105));
	M106: MUX2TO1_1BIT PORT MAP (EM1(106),EM2(106),EMS,SM(106));
	M107: MUX2TO1_1BIT PORT MAP (EM1(107),EM2(107),EMS,SM(107));
	M108: MUX2TO1_1BIT PORT MAP (EM1(108),EM2(108),EMS,SM(108));
	M109: MUX2TO1_1BIT PORT MAP (EM1(109),EM2(109),EMS,SM(109));
	M110: MUX2TO1_1BIT PORT MAP (EM1(110),EM2(110),EMS,SM(110));
	M111: MUX2TO1_1BIT PORT MAP (EM1(111),EM2(111),EMS,SM(111));
	M112: MUX2TO1_1BIT PORT MAP (EM1(112),EM2(112),EMS,SM(112));
	M113: MUX2TO1_1BIT PORT MAP (EM1(113),EM2(113),EMS,SM(113));
	M114: MUX2TO1_1BIT PORT MAP (EM1(114),EM2(114),EMS,SM(114));
	M115: MUX2TO1_1BIT PORT MAP (EM1(115),EM2(115),EMS,SM(115));
	M116: MUX2TO1_1BIT PORT MAP (EM1(116),EM2(116),EMS,SM(116));
	M117: MUX2TO1_1BIT PORT MAP (EM1(117),EM2(117),EMS,SM(117));
	M118: MUX2TO1_1BIT PORT MAP (EM1(118),EM2(118),EMS,SM(118));
	M119: MUX2TO1_1BIT PORT MAP (EM1(119),EM2(119),EMS,SM(119));
	M120: MUX2TO1_1BIT PORT MAP (EM1(120),EM2(120),EMS,SM(120));
	M121: MUX2TO1_1BIT PORT MAP (EM1(121),EM2(121),EMS,SM(121));
	M122: MUX2TO1_1BIT PORT MAP (EM1(122),EM2(122),EMS,SM(122));
	M123: MUX2TO1_1BIT PORT MAP (EM1(123),EM2(123),EMS,SM(123));
	M124: MUX2TO1_1BIT PORT MAP (EM1(124),EM2(124),EMS,SM(124));
	M125: MUX2TO1_1BIT PORT MAP (EM1(125),EM2(125),EMS,SM(125));
	M126: MUX2TO1_1BIT PORT MAP (EM1(126),EM2(126),EMS,SM(126));
	M127: MUX2TO1_1BIT PORT MAP (EM1(127),EM2(127),EMS,SM(127)); 
end MUX2TO1_128BIT;
