library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity SUMADOR2T01_32BITSMOD32 is
	 port(
		 ESA : in STD_LOGIC_VECTOR(31 downto 0);
		 ESB : in STD_LOGIC_VECTOR(31 downto 0);
		 SS : out STD_LOGIC_VECTOR(31 downto 0)
	     );
end SUMADOR2T01_32BITSMOD32;
 
architecture SUMADOR2T01_32BITSMOD32 of SUMADOR2T01_32BITSMOD32 is
signal TSS: STD_LOGIC_VECTOR (32 DOWNTO 0);
begin	
	TSS <= ('0' & ESA) + ('0' & ESB);	 
	 SS <= TSS(31 DOWNTO 0);
end SUMADOR2T01_32BITSMOD32;
