library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity SIGMACHICA0 is
	 port(
		 EX : in  STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SF : out STD_LOGIC_VECTOR(31 DOWNTO 0)
	     );
end SIGMACHICA0;
 
architecture SIGMACHICA0 of SIGMACHICA0 is
COMPONENT XOR2TO1_32BIT is
	 port(
		 EX1 : in STD_LOGIC_VECTOR(31 downto 0);
		 EX2 : in STD_LOGIC_VECTOR(31 downto 0);
		 SX : out STD_LOGIC_VECTOR(31 downto 0)
	     );
end COMPONENT;		   
SIGNAL SX1: STD_LOGIC_VECTOR (31 DOWNTO 0);
begin	   
	XOR1: XOR2TO1_32BIT PORT MAP (
		EX1(31 DOWNTO 25)=>EX( 6 DOWNTO 0),
		EX1(24 DOWNTO  0)=>EX(31 DOWNTO 7),
		EX2(31 DOWNTO 14)=>EX(17 DOWNTO 0),
		EX2(13 DOWNTO  0)=>EX(31 DOWNTO 18),
		SX =>SX1
		);
	XOR2: XOR2TO1_32BIT PORT MAP (
		EX1(31 DOWNTO 29)=>"000",
		EX1(28 DOWNTO  0)=>EX(31 DOWNTO 3),
		EX2=>SX1,
		SX =>SF
		);
end SIGMACHICA0;