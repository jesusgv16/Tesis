library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity SIGMACHICA1 is
	 port(
		 EX : in  STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SF : out STD_LOGIC_VECTOR(31 DOWNTO 0)
	     );
end SIGMACHICA1;
 
architecture SIGMACHICA1 of SIGMACHICA1 is
COMPONENT XOR2TO1_32BIT is
	 port(
		 EX1 : in STD_LOGIC_VECTOR(31 downto 0);
		 EX2 : in STD_LOGIC_VECTOR(31 downto 0);
		 SX : out STD_LOGIC_VECTOR(31 downto 0)
	     );
end COMPONENT;		   
SIGNAL SX1: STD_LOGIC_VECTOR (31 DOWNTO 0);
begin	   
	XOR1: XOR2TO1_32BIT PORT MAP (
		EX1(31 DOWNTO 15)=>EX(16 DOWNTO  0),
		EX1(14 DOWNTO  0)=>EX(31 DOWNTO 17),
		EX2(31 DOWNTO 13)=>EX(18 DOWNTO  0),
		EX2(12 DOWNTO  0)=>EX(31 DOWNTO 19),
		SX =>SX1
		);
	XOR2: XOR2TO1_32BIT PORT MAP (
		EX1(31 DOWNTO 22)=>"0000000000",
		EX1(21 DOWNTO  0)=>EX(31 DOWNTO 10),
		EX2=>SX1,
		SX =>SF
		);
end SIGMACHICA1;