library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity REGTEMP_512BIT is
	 port(
		 ERD : in STD_LOGIC_VECTOR(511 DOWNTO 0);
		 ERW : in STD_LOGIC;
		 CLK : in STD_LOGIC;
		 RST : in STD_LOGIC;
		 SRQ : out STD_LOGIC_VECTOR(511 DOWNTO 0)
	     );
end REGTEMP_512BIT;

architecture REGTEMP_512BIT of REGTEMP_512BIT is
begin
	PROCESS(RST,CLK,ERD,ERW)
	BEGIN		
		IF RST='1' THEN
			SRQ <= x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		ELSIF(RISING_EDGE(CLK)) THEN
			IF (ERW='1') THEN
				SRQ <= ERD;
			END IF;
		END IF;	
	END PROCESS;
end REGTEMP_512BIT;