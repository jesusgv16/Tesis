library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity UnidadProcesamiento is
	 port(
		 WT   : in  STD_LOGIC_VECTOR(31 DOWNTO 0);
		 CLK  : in  STD_LOGIC;
		 RST  : in  STD_LOGIC;	
		 WRB1 : IN  STD_logic ;
		 SELB1: IN  STD_logic ;
		 SELH0: IN  STD_logic ;
		 SELS1: IN  STD_logic ;
		 ADDKT: IN  STd_logic_Vector( 5 DOWNTO  0);
		 HASH : out STD_LOGIC_VECTOR(255 DOWNTO 0)
	     );
end UnidadProcesamiento;

architecture UnidadProcesamiento of UnidadProcesamiento is
COMPONENT MessageSchedule is
	 port(
		 WIN : in  STD_LOGIC_VECTOR(31 downto 0);
		 SEE : in  STD_LOGIC;
		 CLK : in  STD_LOGIC;
		 RST : in  STD_LOGIC;
		 WOU : out STD_LOGIC_VECTOR(31 downto 0)
	     );
end COMPONENT ;
COMPONENT Buffer8x32 is
	 port(
		 H0R : in STD_LOGIC_VECTOR(255 DOWNTO 0);
		 SEL : in STD_LOGIC;
		 ERW : in STD_LOGIC;
		 CLK : in STD_LOGIC;
		 RST : in STD_LOGIC;
		 H0F : out STD_LOGIC_VECTOR(255 DOWNTO 0)
	     );
end COMPONENT;	 
COMPONENT Memory64x32 is
	 port(
		 A : in STD_LOGIC_VECTOR(5 downto 0);
		 SPO : out STD_LOGIC_VECTOR(31 downto 0)
	     );
end COMPONENT;			 
COMPONENT SUMADOR2T01_32BITSMOD32 is
	 port(
		 ESA : in STD_LOGIC_VECTOR(31 downto 0);
		 ESB : in STD_LOGIC_VECTOR(31 downto 0);
		 SS : out STD_LOGIC_VECTOR(31 downto 0)
	     );
end COMPONENT;	 
COMPONENT CH_Function is
	 port(
		 EX : in STD_LOGIC_VECTOR(31 DOWNTO 0);
		 EY : in STD_LOGIC_VECTOR(31 DOWNTO 0);
		 EZ : in STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SF : out STD_LOGIC_VECTOR(31 DOWNTO 0)
	     );
end COMPONENT;		  
COMPONENT MAJ_Function is
	 port(
		 EX : in STD_LOGIC_VECTOR(31 DOWNTO 0);
		 EY : in STD_LOGIC_VECTOR(31 DOWNTO 0);
		 EZ : in STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SF : out STD_LOGIC_VECTOR(31 DOWNTO 0)
	     );
end COMPONENT;
COMPONENT SIGMAGRANDE1 is
	 port(
		 EX : in  STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SF : out STD_LOGIC_VECTOR(31 DOWNTO 0)
	     );
end COMPONENT;		
COMPONENT SIGMAGRANDE0 is
	 port(
		 EX : in  STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SF : out STD_LOGIC_VECTOR(31 DOWNTO 0)
	     );
end COMPONENT;	
COMPONENT REGTEMP_128BIT is
	 port(
		 ERD : in STD_LOGIC_VECTOR(127 downto 0);
		 ERW : in STD_LOGIC;
		 CLK : in STD_LOGIC;
		 RST : in STD_LOGIC;
		 SRQ : out STD_LOGIC_VECTOR(127 downto 0)
	     );
end COMPONENT;
COMPONENT MUX2TO1_128BIT is
	 port(
		 EM1 : in STD_LOGIC_VECTOR(127 downto 0);
		 EM2 : in STD_LOGIC_VECTOR(127 downto 0);
		 EMS : in STD_LOGIC;
		 SM : out STD_LOGIC_VECTOR(127 downto 0)
	     );
end COMPONENT;				   
SIGNAL H0,BUFF,THASH,HASH_O: STD_logic_Vector(255 DOWNTO 0); 
SIGNAL WOUT,KT,SG_1,SG_0,CH,MAJ,SUMHK,SUMWT,SUM1,T1,T2,TE,TA: STD_logic_VEctor (31 DOWNTO 0);
begin					
	MSC: MessageSchedule 	PORT MAP (WT,SELS1,CLK,RST,WOUT);
	BUF: Buffer8x32			PORT MAP (HASH_O,SELB1,WRB1,CLK,RST,H0);
    KTR: Memory64x32		PORT MAP (ADDKT,KT);
	SHK: SUMADOR2T01_32BITSMOD32 PORT MAP (BUFF(255 DOWNTO 224),KT,SUMHK);
	SUW: SUMADOR2T01_32BITSMOD32 PORT MAP (SUMHK,WOUT,SUMWT);
	CHF: CH_Function		PORT MAP (BUFF(159 DOWNTO 128),BUFF(191 DOWNTO 160),BUFF(223 DOWNTO 192),CH);
	SG1: SIGMAGRANDE1		PORT MAP (BUFF(159 DOWNTO 128),SG_1);										 
	SU1: SUMADOR2T01_32BITSMOD32 PORT MAP (CH ,SG_1,SUM1);
	MAF: MAJ_Function		PORT MAP (BUFF( 31 DOWNTO   0),BUFF( 63 DOWNTO  32),BUFF( 95 DOWNTO  64),MAJ);
	SG0: SIGMAGRANDE0		PORT MAP (BUFF( 31 DOWNTO   0),SG_0);
	SU2: SUMADOR2T01_32BITSMOD32 PORT MAP (MAJ,SG_0,T2);
	S1W: SUMADOR2T01_32BITSMOD32 PORT MAP (SUM1,SUMWT,T1);   
	SUE: SUMADOR2T01_32BITSMOD32 PORT MAP (T1,BUFF(127 DOWNTO 96),TE);
	SUA: SUMADOR2T01_32BITSMOD32 PORT MAP (T1,T2,TA);	 
	RH1: REGTEMP_128BIT 	PORT MAP (
		ERD(127 DOWNTO  96) => BUFF(223 DOWNTO 192),
		ERD( 95 DOWNTO  64) => BUFF(191 DOWNTO 160),
		ERD( 63 DOWNTO  32) => BUFF(159 DOWNTO 128),
		ERD( 31 DOWNTO   0) => TE,
		ERW => '1',
		CLK => CLK,
		RST => RST,
		SRQ => THASH(255 DOWNTO 128));
	RH2: REGTEMP_128BIT		PORT MAP (
     	ERD(127 DOWNTO  96) => BUFF( 95 DOWNTO  64),
		ERD( 95 DOWNTO  64) => BUFF( 63 DOWNTO  32),
		ERD( 63 DOWNTO  32) => BUFF( 31 DOWNTO   0),
		ERD( 31 DOWNTO   0) => TA,
		ERW => '1',
		CLK => CLK,
		RST => RST,
		SRQ => THASH(127 DOWNTO   0));					 
	MU1: MUX2TO1_128BIT	PORT MAP (THASH(255 DOWNTO 128),H0(255 DOWNTO 128),SELH0,BUFF(255 DOWNTO 128));
	MU2: MUX2TO1_128BIT PORT MAP (THASH(127 DOWNTO   0),H0(127 DOWNTO   0),SELH0,BUFF(127 DOWNTO   0));
	
	HA1: SUMADOR2T01_32BITSMOD32 PORT MAP (BUFF(255 DOWNTO 224),THASH(255 DOWNTO 224),HASH_O(255 DOWNTO 224));
	HA2: SUMADOR2T01_32BITSMOD32 PORT MAP (BUFF(223 DOWNTO 192),THASH(223 DOWNTO 192),HASH_O(223 DOWNTO 192));
	HA3: SUMADOR2T01_32BITSMOD32 PORT MAP (BUFF(191 DOWNTO 160),THASH(191 DOWNTO 160),HASH_O(191 DOWNTO 160));
	HA4: SUMADOR2T01_32BITSMOD32 PORT MAP (BUFF(159 DOWNTO 128),THASH(159 DOWNTO 128),HASH_O(159 DOWNTO 128));
	HA5: SUMADOR2T01_32BITSMOD32 PORT MAP (BUFF(127 DOWNTO  96),THASH(127 DOWNTO  96),HASH_O(127 DOWNTO  96));
	HA6: SUMADOR2T01_32BITSMOD32 PORT MAP (BUFF( 95 DOWNTO  64),THASH( 95 DOWNTO  64),HASH_O( 95 DOWNTO  64));
	HA7: SUMADOR2T01_32BITSMOD32 PORT MAP (BUFF( 63 DOWNTO  32),THASH( 63 DOWNTO  32),HASH_O( 63 DOWNTO  32));
	HA8: SUMADOR2T01_32BITSMOD32 PORT MAP (BUFF( 31 DOWNTO   0),THASH( 31 DOWNTO   0),HASH_O( 31 DOWNTO   0));
	HASH <= HASH_O;
end UnidadProcesamiento;